`timescale 1ns / 1ps

module drone_top_tb;

    reg clk;
    reg rst_n;
    reg RxD;
    reg signal_INT;
    wire scl;
    wire sda;           // ��Ϊ wire���� I?C ���豸����
    wire pwm_1, pwm_2, pwm_3, pwm_4;

    // ģ�� I?C �豸���� sda������ MPU6050��
    reg sda_drive = 1;  // Ĭ�ϸߵ�ƽ���ͷţ�
    reg sda_dir = 0;    // 0: �ͷţ�����̬����1: ����
    assign sda = sda_dir ? sda_drive : 1'bz;  // ��̬����
    //assign sda = sda_dir ? sda_drive : 1'b1;  // ��̬����,����ʱ������ȫ1����

    // ʵ��������ģ��
    drone_top uut (
        .clk(clk),
        .rst_n(rst_n),
        .scl(scl),
        .sda(sda),
        .signal_INT(signal_INT),
        .pwm_1(pwm_1),
        .pwm_2(pwm_2),
        .pwm_3(pwm_3),
        .pwm_4(pwm_4),
        .RxD(RxD) 
    );

    // ����ʱ��
    always #10 clk = ~clk;

    // ģ�⴮������
    task send_uart_byte(input [7:0] data);
        integer i;
        begin
            RxD = 0; // ��ʼλ
            #8680;  // 115200 baud -> һ��bitʱ��Լ8.68us
            for (i = 0; i < 8; i = i + 1) begin
                RxD = data[i];
                #8680;
            end
            RxD = 1; // ֹͣλ
            #8680;
        end
    endtask

    // ���Թ���
    initial begin
        clk = 0;
        rst_n = 0;
        RxD = 1;
        sda_dir = 0;  // ��ʼ�ͷ� sda

        // ��λ
        #50 rst_n = 1;

        #100 signal_INT = 1;

        // ���ʹ��������� 8'h01��
        #1000 send_uart_byte(8'h0A); // START_BYTE
        #1000 send_uart_byte(8'h04); // ǰ��
        #1000 send_uart_byte(8'h08); // STOP_BYTE

        #100000 signal_INT = 0;
        #500000 signal_INT = 1;
        #100000 signal_INT = 0;

        #500000 signal_INT = 1;
        #100000 signal_INT = 0;

        // ��������һ��ʱ��
        #100000;
        
        // ֹͣ����
        $finish;
    end
endmodule